`timescale 1ns / 1ps

module core_sim;
    reg clk, rst;

    RV32core core(
        .clk(clk),
        .rst(rst)
    );

    initial begin
        clk = 0;
        rst = 1;
        #2 rst = 0;
    end
    always #1 clk = ~clk;

    // Signals to probe

    wire [31:0] PC_IF, inst_IF, PC_ID, inst_ID, PC_EXE, inst_EXE, PC_WB, inst_WB;

    assign PC_IF    = core.PC_IF;
    assign inst_IF  = core.inst_IF;
    assign PC_ID    = core.PC_ID;
    assign inst_ID  = core.inst_ID;
    assign PC_EXE   = core.PC_EXE;
    assign inst_EXE = core.inst_EXE;
    assign PC_WB    = core.PC_WB;
    assign inst_WB  = core.inst_WB;

    wire branch, JALR, regWrite_ID, memWrite_ID, MIO_ID, ALUSrc_A_ID, ALUSrc_B_ID, dataToReg_ID;
    
    // x1~x31
    wire [31:0] reg_x [1:31];

    assign branch       = core.branch;
    assign JALR         = core.ID_stage.JALR;
    assign regWrite_ID  = core.regWrite_ID;
    assign memWrite_ID  = core.memWrite_ID;
    assign MIO_ID       = core.MIO_ID;
    assign ALUSrc_A_ID  = core.ALUSrc_A_ID;
    assign ALUSrc_B_ID  = core.ALUSrc_B_ID;
    assign dataToReg_ID = core.dataToReg_ID;
    genvar i;
    generate
        for (i=1; i<32; i=i+1) begin
            assign reg_x[i] = core.ID_stage.register.register[i];
        end
    endgenerate

    // Check results

    integer pass;

    initial begin
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000000 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000000 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000000 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000000 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000000 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000000 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000000 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000000 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000004 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00402103 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000000 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000000 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000008 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00802203 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000004 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00402103 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000000 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000000c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x004100b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000008 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00802203 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000004 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00402103 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000010 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xfff08093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000000c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x004100b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000008 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00802203 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000010 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xfff08093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000000c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x004100b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000000c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000000 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000014) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000014 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00c02283) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00c02283 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000010 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_ID expected 0xfff08093 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000000c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x004100b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000004 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00402103 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000000 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000018) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000018 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01002303) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01002303 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000014) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000014 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00c02283) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00c02283 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000010 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0xfff08093 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000008 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00802203 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000001c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000001c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01402383) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01402383 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000018) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000018 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01002303) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01002303 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000014) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000014 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00c02283) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00c02283 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000000c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000020) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000020 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h402200b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x402200b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000001c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000001c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01402383) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01402383 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000018) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000018 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01002303) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01002303 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000000c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x004100b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000018) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000018 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000024) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000024 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h002220b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x002220b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000020) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000020 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h402200b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x402200b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000001c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000001c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01402383) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01402383 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000010 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_WB expected 0xfff08093 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000017) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000017 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000000 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000028) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000028 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h004120b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x004120b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000024) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000024 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h002220b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x002220b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000020) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000020 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h402200b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x402200b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000014) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000014 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00c02283) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00c02283 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000017) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000017 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x00000000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000002c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000002c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h4023d0b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x4023d0b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000028) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000028 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h004120b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x004120b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000024) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000024 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h002220b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x002220b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000018) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000018 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01002303) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01002303 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000017) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000017 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000030) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000030 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h007330b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x007330b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000002c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000002c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h4023d0b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x4023d0b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000028) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000028 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h004120b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x004120b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000001c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000001c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01402383) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01402383 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000017) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000017 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000034) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000034 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hffd38093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xffd38093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000030) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000030 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h007330b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x007330b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000002c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000002c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h4023d0b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x4023d0b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000020) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000020 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h402200b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x402200b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000008 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000038) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000038 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00f22093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00f22093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000034) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000034 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'hffd38093) begin pass = 0; $display("Time: %3dns, inst_ID expected 0xffd38093 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000030) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000030 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h007330b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x007330b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000024) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000024 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h002220b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x002220b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000003c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000003c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00225093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00225093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000038) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000038 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00f22093) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00f22093 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000034) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000034 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'hffd38093) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0xffd38093 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000028) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000028 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h004120b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x004120b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000001) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000001 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000040) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000040 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h40c35093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x40c35093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000003c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000003c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00225093) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00225093 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000038) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000038 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00f22093) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00f22093 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000002c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000002c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h4023d0b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x4023d0b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000044) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000044 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01802403) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01802403 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000040) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000040 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h40c35093) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x40c35093 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000003c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000003c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00225093) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00225093 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000030) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000030 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h007330b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x007330b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000048 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00802e23) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00802e23 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000044) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000044 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01802403) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01802403 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000040) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000040 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h40c35093) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x40c35093 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000034) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000034 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'hffd38093) begin pass = 0; $display("Time: %3dns, inst_WB expected 0xffd38093 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hfffffffd) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xfffffffd but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000004c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000004c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01c02083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01c02083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000048 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00802e23) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00802e23 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000044) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000044 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01802403) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01802403 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000038) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000038 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00f22093) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00f22093 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000000 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000004c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000004c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01c02083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01c02083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000048 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00802e23) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00802e23 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000048 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000003c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000003c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00225093) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00225093 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000004) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000004 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000050) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000050 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h02801023) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x02801023 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000004c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000004c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01c02083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01c02083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000048 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00802e23) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00802e23 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000040) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000040 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h40c35093) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x40c35093 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hfffffff0) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xfffffff0 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x00000000 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000054) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000054 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h02002083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x02002083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000050) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000050 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h02801023) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x02801023 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000004c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000004c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01c02083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01c02083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000044) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000044 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01802403) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01802403 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hfffffff0) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xfffffff0 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000058) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000058 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h02800223) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x02800223 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000054) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000054 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h02002083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x02002083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000050) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000050 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h02801023) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x02801023 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000048 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hfffffff0) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xfffffff0 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000005c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000005c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h02402083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x02402083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000058) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000058 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h02800223) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x02800223 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000054) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000054 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h02002083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x02002083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000048) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000048 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00802e23) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00802e23 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hfffffff0) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xfffffff0 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000060) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000060 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01a01083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01a01083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000005c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000005c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h02402083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x02402083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000058) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000058 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h02800223) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x02800223 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000004c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000004c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01c02083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01c02083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000f0f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000f0f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000064) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000064 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01a05083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01a05083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000060) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000060 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01a01083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01a01083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000005c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000005c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h02402083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x02402083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000050) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000050 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h02801023) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x02801023 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000f0f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000f0f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000068) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000068 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01b00083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01b00083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000064) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000064 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01a05083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01a05083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000060) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000060 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01a01083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01a01083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000054) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000054 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h02002083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x02002083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000006c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000006c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h01b04083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x01b04083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000068) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000068 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01b00083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01b00083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000064) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000064 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01a05083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01a05083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000058) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000058 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h02800223) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x02800223 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000070) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000070 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hffff0097) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xffff0097 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000006c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000006c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h01b04083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x01b04083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000068) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000068 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01b00083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01b00083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000005c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000005c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h02402083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x02402083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000074) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000074 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000070) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000070 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'hffff0097) begin pass = 0; $display("Time: %3dns, inst_ID expected 0xffff0097 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000006c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000006c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h01b04083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x01b04083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000060) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000060 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01a01083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01a01083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h00000f0f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x00000f0f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000078) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000078 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000074) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000074 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000070) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000070 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'hffff0097) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0xffff0097 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000064) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000064 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01a05083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01a05083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000007c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000007c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000078) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000078 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000074) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000074 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000068) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000068 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01b00083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01b00083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000080) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000080 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h02c02083) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x02c02083 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000007c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000007c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000078) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000078 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000006c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000006c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h01b04083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x01b04083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h0000000f) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x0000000f but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000084) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000084 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03802103) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03802103 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000080) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000080 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h02c02083) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x02c02083 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000007c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000007c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000070) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000070 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'hffff0097) begin pass = 0; $display("Time: %3dns, inst_WB expected 0xffff0097 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hffff0070) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xffff0070 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000088 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h002081ab) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x002081ab but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000084) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000084 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h03802103) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x03802103 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000080) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000080 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h02c02083) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x02c02083 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000074) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000074 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hffff0070) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xffff0070 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000008c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000008c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03002203) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03002203 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000088 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h002081ab) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x002081ab but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000084) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000084 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h03802103) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x03802103 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000078) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000078 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hffff0070) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xffff0070 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000008c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000008c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03002203) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03002203 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000088 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h002081ab) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x002081ab but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000088 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000007c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000007c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'hffff0070) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0xffff0070 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000090) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000090 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03c02283) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03c02283 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000008c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000008c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h03002203) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x03002203 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000088 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h002081ab) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x002081ab but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000080) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000080 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h02c02083) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x02c02083 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h00000008) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x00000008 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000094 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h0052032b) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x0052032b but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000090) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000090 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h03c02283) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x03c02283 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000008c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000008c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h03002203) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x03002203 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000084) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000084 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h03802103) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x03802103 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000098) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000098 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03402383) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03402383 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000094 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h0052032b) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x0052032b but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000090) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000090 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h03c02283) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x03c02283 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000088 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00000000 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000098) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000098 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h03402383) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x03402383 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000094 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h0052032b) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x0052032b but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000094 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000088) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000088 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h002081ab) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x002081ab but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h00000010) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x00000010 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000009c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000009c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h04002403) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x04002403 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000098) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000098 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h03402383) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x03402383 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000094 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h0052032b) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x0052032b but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000008c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000008c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h03002203) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x03002203 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h00000014) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x00000014 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000a0 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h008384ab) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x008384ab but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000009c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000009c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h04002403) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x04002403 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000098) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000098 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h03402383) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x03402383 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000090) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000090 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h03c02283) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x03c02283 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000a4) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000a4 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h006181b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x006181b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000a0 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h008384ab) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x008384ab but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000009c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000009c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h04002403) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x04002403 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000094 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'hffff0000) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0xffff0000 but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000a4) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000a4 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h006181b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x006181b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000a0 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h008384ab) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x008384ab but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000a0 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000094) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000094 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h0052032b) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x0052032b but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x00000000 but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000a8 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h009181b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x009181b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000a4) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000a4 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h006181b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x006181b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000a0 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h008384ab) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x008384ab but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000098) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000098 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h03402383) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x03402383 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'hff000f0f) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0xff000f0f but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000ac) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000ac but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h04302223) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x04302223 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000a8 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h009181b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x009181b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000a4) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000a4 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h006181b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x006181b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h0000009c) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x0000009c but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h04002403) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x04002403 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000ac) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000ac but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h04302223) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x04302223 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000a8 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h009181b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x009181b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000a8 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000a0 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00000000 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000b0) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000b0 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000ac) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000ac but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h04302223) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x04302223 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000a8 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h009181b3) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x009181b3 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000a0) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000a0 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h008384ab) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x008384ab but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000093b) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000093b but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000b4) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000b4 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000b0) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000b0 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000ac) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000ac but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h04302223) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x04302223 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000a4) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000a4 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h006181b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x006181b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00006138) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00006138 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000b8) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000b8 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000b4) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000b4 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000b0) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000b0 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000a8 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000000 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h00006138) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x00006138 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000bc but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hf45ff06f) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xf45ff06f but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000b8) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000b8 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000b4) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000b4 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000a8) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000a8 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h009181b3) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x009181b3 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h000000c0) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x000000c0 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hxxxxxxxx) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xxxxxxxxx but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000bc but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'hf45ff06f) begin pass = 0; $display("Time: %3dns, inst_ID expected 0xf45ff06f but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000b8) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000b8 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000ac) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000ac but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h04302223) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x04302223 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000000 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00000013 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x000000bc but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000bc but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'hf45ff06f) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0xf45ff06f but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000b0) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000b0 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000004 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00402103 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000000 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00000013 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x000000bc but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000b4) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000b4 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000008 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x00802203 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000004 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00402103 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000000 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000013 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000b8) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000b8 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x0000000c but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_IF expected 0x004100b3 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x00000008 but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x00802203 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000004) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000004 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00402103) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00402103 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000bc but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'hf45ff06f) begin pass = 0; $display("Time: %3dns, inst_WB expected 0xf45ff06f but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000010 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xfff08093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000000c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x004100b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h00000008) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x00000008 but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00802203) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00802203 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h000000bc) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x000000bc but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        pass = 1;
        if (PC_IF !== 32'h00000010) begin pass = 0; $display("Time: %3dns, PC_IF expected 0x00000010 but get 0x%08x", $time, PC_IF); end
        if (inst_IF !== 32'hfff08093) begin pass = 0; $display("Time: %3dns, inst_IF expected 0xfff08093 but get 0x%08x", $time, inst_IF); end
        if (PC_ID !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_ID expected 0x0000000c but get 0x%08x", $time, PC_ID); end
        if (inst_ID !== 32'h004100b3) begin pass = 0; $display("Time: %3dns, inst_ID expected 0x004100b3 but get 0x%08x", $time, inst_ID); end
        if (PC_EXE !== 32'h0000000c) begin pass = 0; $display("Time: %3dns, PC_EXE expected 0x0000000c but get 0x%08x", $time, PC_EXE); end
        if (inst_EXE !== 32'h00000000) begin pass = 0; $display("Time: %3dns, inst_EXE expected 0x00000000 but get 0x%08x", $time, inst_EXE); end
        if (PC_WB !== 32'h00000000) begin pass = 0; $display("Time: %3dns, PC_WB expected 0x00000000 but get 0x%08x", $time, PC_WB); end
        if (inst_WB !== 32'h00000013) begin pass = 0; $display("Time: %3dns, inst_WB expected 0x00000013 but get 0x%08x", $time, inst_WB); end
        if (reg_x[1] !== 32'h11223344) begin pass = 0; $display("Time: %3dns, reg_x[1] expected 0x11223344 but get 0x%08x", $time, reg_x[1]); end
        if (reg_x[2] !== 32'h20250306) begin pass = 0; $display("Time: %3dns, reg_x[2] expected 0x20250306 but get 0x%08x", $time, reg_x[2]); end
        if (reg_x[3] !== 32'h0000f581) begin pass = 0; $display("Time: %3dns, reg_x[3] expected 0x0000f581 but get 0x%08x", $time, reg_x[3]); end
        if (reg_x[4] !== 32'h55667788) begin pass = 0; $display("Time: %3dns, reg_x[4] expected 0x55667788 but get 0x%08x", $time, reg_x[4]); end
        if (reg_x[5] !== 32'h18970521) begin pass = 0; $display("Time: %3dns, reg_x[5] expected 0x18970521 but get 0x%08x", $time, reg_x[5]); end
        if (reg_x[6] !== 32'h000057fd) begin pass = 0; $display("Time: %3dns, reg_x[6] expected 0x000057fd but get 0x%08x", $time, reg_x[6]); end
        if (reg_x[7] !== 32'h99aabbcc) begin pass = 0; $display("Time: %3dns, reg_x[7] expected 0x99aabbcc but get 0x%08x", $time, reg_x[7]); end
        if (reg_x[8] !== 32'h21121480) begin pass = 0; $display("Time: %3dns, reg_x[8] expected 0x21121480 but get 0x%08x", $time, reg_x[8]); end
        if (reg_x[9] !== 32'h00009449) begin pass = 0; $display("Time: %3dns, reg_x[9] expected 0x00009449 but get 0x%08x", $time, reg_x[9]); end
        if (reg_x[10] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[10] expected 0x00000000 but get 0x%08x", $time, reg_x[10]); end
        if (reg_x[11] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[11] expected 0x00000000 but get 0x%08x", $time, reg_x[11]); end
        if (reg_x[12] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[12] expected 0x00000000 but get 0x%08x", $time, reg_x[12]); end
        if (reg_x[13] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[13] expected 0x00000000 but get 0x%08x", $time, reg_x[13]); end
        if (reg_x[14] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[14] expected 0x00000000 but get 0x%08x", $time, reg_x[14]); end
        if (reg_x[15] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[15] expected 0x00000000 but get 0x%08x", $time, reg_x[15]); end
        if (reg_x[16] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[16] expected 0x00000000 but get 0x%08x", $time, reg_x[16]); end
        if (reg_x[17] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[17] expected 0x00000000 but get 0x%08x", $time, reg_x[17]); end
        if (reg_x[18] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[18] expected 0x00000000 but get 0x%08x", $time, reg_x[18]); end
        if (reg_x[19] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[19] expected 0x00000000 but get 0x%08x", $time, reg_x[19]); end
        if (reg_x[20] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[20] expected 0x00000000 but get 0x%08x", $time, reg_x[20]); end
        if (reg_x[21] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[21] expected 0x00000000 but get 0x%08x", $time, reg_x[21]); end
        if (reg_x[22] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[22] expected 0x00000000 but get 0x%08x", $time, reg_x[22]); end
        if (reg_x[23] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[23] expected 0x00000000 but get 0x%08x", $time, reg_x[23]); end
        if (reg_x[24] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[24] expected 0x00000000 but get 0x%08x", $time, reg_x[24]); end
        if (reg_x[25] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[25] expected 0x00000000 but get 0x%08x", $time, reg_x[25]); end
        if (reg_x[26] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[26] expected 0x00000000 but get 0x%08x", $time, reg_x[26]); end
        if (reg_x[27] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[27] expected 0x00000000 but get 0x%08x", $time, reg_x[27]); end
        if (reg_x[28] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[28] expected 0x00000000 but get 0x%08x", $time, reg_x[28]); end
        if (reg_x[29] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[29] expected 0x00000000 but get 0x%08x", $time, reg_x[29]); end
        if (reg_x[30] !== 32'h00000000) begin pass = 0; $display("Time: %3dns, reg_x[30] expected 0x00000000 but get 0x%08x", $time, reg_x[30]); end
        if (reg_x[31] !== 32'h0000000) begin pass = 0; $display("Time: %3dns, reg_x[31] expected 0x0000000 but get 0x%08x", $time, reg_x[31]); end
        if (pass == 1) begin $display("Time: %3dns, pass.", $time); end else begin @(posedge clk); $stop(); end
        @(posedge clk);
        $display("All samples passed! Congrats!");
        $stop();
    end

endmodule