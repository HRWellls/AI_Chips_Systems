` timescale 1ns / 1ps

module Vdot(
    input clk,                                        
    input rst,
    input EN,                                           
    input[31:0] A, B,
    output[31:0] res
);

// [Topic 1] Please finish the code of vector dot product that requires 3 cycles for execution.
// You can use the Mult4 module in common/MULT4.v to implement the multiplication of 4-bit numbers.

// You may add some code here...

assign res = // Complete the signal here.

endmodule